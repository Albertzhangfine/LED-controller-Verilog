module ledd(clk,rst,led,state_ctrl);  
  
input clk ;  
input rst ;  
input state_ctrl;
output reg [15:0]led ;  
  
reg[5:0] state;  
reg[3:0] state_k;

always @ ( posedge clk or negedge rst or negedge state_ctrl)
begin

	if(!rst)
		begin
			led<=16'b1111111111111111;
			state<=0;
		end
	else 
	begin
	  if(!state_ctrl)
	     begin
			led<=16'b0000000000000000;
			state<=0;
			
		  end
	  else
	   begin
		case (state_k)
			0:begin
			case(state)
				0:begin
					led<='b0111111111111111;
					state<=1;
				end
				1:begin
					led<='b1011111111111111;
					state<=2;	
				end
				2:begin
					led<='b1101111111111111;	
					state<=3;			
				end
				3:begin
					led<='b1110111111111111;
					state<=4;	
				end
				4:begin
					led<='b1111011111111111;
					state<=5;
					end
				5:begin
					led<='b1111101111111111;
					state<=6;
					end
				6:begin
					led<='b1111110111111111;
					state<=7;
					end
				7:begin
					led<='b1111111011111111;
					state<=8;
					end
				8:begin
					led<='b1111111101111111;
					state<=9;
					end
				9:begin
					led<='b1111111110111111;
					state<=10;
					end
				10:begin
					led<='b1111111111011111;
					state<=11;
					end
				11:begin
					led<='b1111111111101111;
					state<=12;
					end
				12:begin
					led<='b1111111111110111;
					state<=13;
					end
				13:begin
					led<='b1111111111111011;
					state<=14;
					end
				14:begin
					led<='b1111111111111101;
					state<=15;
					end
				15:begin
					led<='b1111111111111110;
					state<=16;
					end
				default: 
					state<=0;
				endcase
				state_k<=1;
			end
			1:begin
			case(state)
				0:begin
					led<='b0111111111111110;
					state<=1;
				end
				1:begin
					led<='b1011111111111101;
					state<=2;	
				end
				2:begin
					led<='b1101111111111011;	
					state<=3;			
				end
				3:begin
					led<='b1110111111110111;
					state<=4;	
				end
				4:begin
					led<='b1111011111101111;
					state<=5;
					end
				5:begin
					led<='b1111101111011111;
					state<=6;
					end
				6:begin
					led<='b1111110110111111;
					state<=7;
					end
				7:begin
					led<='b1111111001111111;
					state<=8;
					end
				
				default: 
					state<=0;
				endcase
				state_k<=2;
			
			end
			2:begin
			case(state)
				0:begin
					led<='b0011111111111100;
					state<=1;
				end
				1:begin
					led<='b1001111111111001;
					state<=2;	
				end
				2:begin
					led<='b1100111111110011;	
					state<=3;			
				end
				3:begin
					led<='b1110011111100111;
					state<=4;	
				end
				4:begin
					led<='b1111001111001111;
					state<=5;
					end
				5:begin
					led<='b1111100110011111;
					state<=6;
					end
				6:begin
					led<='b1111110000111111;
					state<=7;
					end
				7:begin
					led<='b1111111001111111;
					state<=8;
					end
				
				default: 
					state<=0;
				endcase
				state_k<=3;
			end
			3:begin
			case(state)
				0:begin
					led<='b0111111111111111;
					state<=1;
				end
				1:begin
					led<='b1011111111111111;
					state<=2;	
				end
				2:begin
					led<='b1101111111111111;	
					state<=3;			
				end
				3:begin
					led<='b1110111111111111;
					state<=4;	
				end
				4:begin
					led<='b1111011111111111;
					state<=5;
					end
				5:begin
					led<='b1111101111111111;
					state<=6;
					end
				6:begin
					led<='b1111110111111111;
					state<=7;
					end
				7:begin
					led<='b1111111011111111;
					state<=8;
					end
				8:begin
					led<='b1111111101111111;
					state<=9;
					end
				9:begin
					led<='b1111111110111111;
					state<=10;
					end
				10:begin
					led<='b1111111111011111;
					state<=11;
					end
				11:begin
					led<='b1111111111101111;
					state<=12;
					end
				12:begin
					led<='b1111111111110111;
					state<=13;
					end
				13:begin
					led<='b1111111111111011;
					state<=14;
					end
				14:begin
					led<='b1111111111111101;
					state<=15;
					end
				15:begin
					led<='b1111111111111110;
					state<=16;
					end
				default: 
					state<=0;
				endcase
				state_k<=4;
			end
			4:begin
			case(state)
				0:begin
					led<='b0111111111111111;
					state<=1;
				end
				1:begin
					led<='b1011111111111111;
					state<=2;	
				end
				2:begin
					led<='b1101111111111111;	
					state<=3;			
				end
				3:begin
					led<='b1110111111111111;
					state<=4;	
				end
				4:begin
					led<='b1111011111111111;
					state<=5;
					end
				5:begin
					led<='b1111101111111111;
					state<=6;
					end
				6:begin
					led<='b1111110111111111;
					state<=7;
					end
				7:begin
					led<='b1111111011111111;
					state<=8;
					end
				8:begin
					led<='b1111111101111111;
					state<=9;
					end
				9:begin
					led<='b1111111110111111;
					state<=10;
					end
				10:begin
					led<='b1111111111011111;
					state<=11;
					end
				11:begin
					led<='b1111111111101111;
					state<=12;
					end
				12:begin
					led<='b1111111111110111;
					state<=13;
					end
				13:begin
					led<='b1111111111111011;
					state<=14;
					end
				14:begin
					led<='b1111111111111101;
					state<=15;
					end
				15:begin
					led<='b1111111111111110;
					state<=16;
					end
				default: 
					state<=0;
				endcase
				state_k<=5;
			end
			5:begin
			case(state)
				0:begin
					led<='b0111111111111111;
					state<=1;
				end
				1:begin
					led<='b1011111111111111;
					state<=2;	
				end
				2:begin
					led<='b1101111111111111;	
					state<=3;			
				end
				3:begin
					led<='b1110111111111111;
					state<=4;	
				end
				4:begin
					led<='b1111011111111111;
					state<=5;
					end
				5:begin
					led<='b1111101111111111;
					state<=6;
					end
				6:begin
					led<='b1111110111111111;
					state<=7;
					end
				7:begin
					led<='b1111111011111111;
					state<=8;
					end
				8:begin
					led<='b1111111101111111;
					state<=9;
					end
				9:begin
					led<='b1111111110111111;
					state<=10;
					end
				10:begin
					led<='b1111111111011111;
					state<=11;
					end
				11:begin
					led<='b1111111111101111;
					state<=12;
					end
				12:begin
					led<='b1111111111110111;
					state<=13;
					end
				13:begin
					led<='b1111111111111011;
					state<=14;
					end
				14:begin
					led<='b1111111111111101;
					state<=15;
					end
				15:begin
					led<='b1111111111111110;
					state<=16;
					end
				default: 
					state<=0;
				endcase
				state_k<=0;
			end
			default: 
					state_k<=0;
			endcase
			
	   end
	end
end
endmodule  
