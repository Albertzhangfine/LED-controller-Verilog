module led_16(clk,rst,speed,state_ctrl,led,clk_show);

input clk ;
input rst ;
input speed ;//速度控制，0为快节奏，1为慢节奏
input state_ctrl ;//花色控制，1为花色循环变化，0为花色不变,高有效
output reg [15:0] led ;

reg [5:0] state ;
reg [15:0] counter ;
output reg clk_show;

always @ ( posedge clk or negedge rst or negedge speed)
begin
	if(!rst)
		begin
			clk_show<=0;
			counter<=0;
		end
	case(speed)
	  0:begin
	    	if(counter<10)
		    	counter<=counter+1;
		   else
			begin
				counter<=0;			
				clk_show<=~clk_show;
			end
	  end
	 1:begin 
	      if(counter<40)
		    	counter<=counter+1;
		   else
			begin
				counter<=0;			
				clk_show<=~clk_show;
			end
     end
	 endcase
end
always @ ( posedge clk_show or negedge rst or negedge state_ctrl)
begin

	if(!rst)
		begin
			led<=16'b1111111111111111;
			state<=0;
		end
	else 
	begin
	  if(!state_ctrl)
	     begin
			led<=16'b0000000000000000;
			state<=0;
			
		  end
	  else
	   begin
		case(state)
		//1
			0:begin
				led<='b0111111111111111;
				state<=1;
			end
			1:begin
				led<='b1011111111111111;
				state<=2;	
			end
			2:begin
				led<='b1101111111111111;	
				state<=3;			
			end
			3:begin
				led<='b1110111111111111;
				state<=4;	
			end
			4:begin
				led<='b1111011111111111;
				state<=5;
				end
			5:begin
				led<='b1111101111111111;
				state<=6;
				end
			6:begin
				led<='b1111110111111111;
				state<=7;
				end
			7:begin
				led<='b1111111011111111;
				state<=8;
				end
			8:begin
				led<='b1111111101111111;
				state<=9;
				end
			9:begin
				led<='b1111111110111111;
				state<=10;
				end
			10:begin
				led<='b1111111111011111;
				state<=11;
				end
			11:begin
				led<='b1111111111101111;
				state<=12;
				end
			12:begin
				led<='b1111111111110111;
				state<=13;
				end
			13:begin
				led<='b1111111111111011;
				state<=14;
				end
			14:begin
				led<='b1111111111111101;
				state<=15;
				end
			15:begin
				led<='b1111111111111110;
				state<=16;
				end
				//2
			16:begin
				led<='b0111111111111110;
				state<=17;
			end
			17:begin
				led<='b1011111111111101;
				state<=18;	
			end
			18:begin
				led<='b1101111111111011;	
				state<=19;			
			end
			19:begin
				led<='b1110111111110111;
				state<=20;	
			end
			20:begin
				led<='b1111011111101111;
				state<=21;
				end
			21:begin
				led<='b1111101111011111;
				state<=22;
				end
			22:begin
				led<='b1111110110111111;
				state<=23;
				end
			23:begin
				led<='b1111111001111111;
				state<=24;
				end
				//3
			24:begin
				led<='b0011111111111100;
				state<=25;
			end
			25:begin
				led<='b1001111111111001;
				state<=26;	
			end
			26:begin
				led<='b1100111111110011;	
				state<=27;			
			end
			27:begin
				led<='b1110011111100111;
				state<=28;	
			end
			28:begin
				led<='b1111001111001111;
				state<=29;
				end
			29:begin
				led<='b1111100110011111;
				state<=30;
				end
			30:begin
				led<='b1111110000111111;
				state<=31;
				end
			31:begin
				led<='b1111111001111111;
				state<=0;
				end
				//4
			32:begin
				led<='b0111111111111111;
				state<=33;
				end
			33:begin
				led<='b1111111111111101;
				state<=34;
				end
			34:begin
				led<='b1101111111111111;
				state<=35;
				end
			35:begin
				led<='b1111111111110111;
				state<=36;
				end
			36:begin
				led<='b1111011111111111;
				state<=37;
				end
			37:begin
				led<='b1111111110111111;
				state<=38;
				end
			38:begin
				led<='b1111110111111111;
				state<=39;
				end
			39:begin
				led<='b1111111011111111;
				state<=40;
				end
				//5
			40:begin
				led<='b1111111001111111;
				state<=41;
				end
			41:begin
				led<='b1111110110111111;
				state<=42;
				end
			42:begin
				led<='b1111101111011111;
				state<=43;
				end
			43:begin
				led<='b1111011111101111;
				state<=44;
				end
			44:begin
				led<='b1110111111110111;
				state<=45;
				end
			45:begin
				led<='b1101111111111011;
				state<=46;
				end
			46:begin
				led<='b1011111111111101;
				state<=47;
				end
			47:begin
				led<='b0111111111111110;
				state<=48;
				end
				//6
			48:begin
				led<='b1111111001111111;
				state<=49;
				end
			49:begin
				led<='b1111110110111111;
				state<=50;
				end
			50:begin
				led<='b1111101111011111;
				state<=51;
				end
			51:begin
				led<='b1111011111101111;
				state<=52;
				end
			52:begin
				led<='b1110111111110111;
				state<=53;
				end
			53:begin
				led<='b1101111111111011;
				state<=54;
				end
			54:begin
				led<='b1011111111111101;
				state<=55;
				end
			55:begin
				led<='b0111111111111110;
				state<=0;
				end
			
			default: 
				state<=0;
			endcase
			
	   end
	end
end
endmodule

